// +FHDR----------------------------------------------------------------------------
//                 Copyright (c) 2022 
//                       ALL RIGHTS RESERVED
// ---------------------------------------------------------------------------------
// Filename      : ysyx_22041752_ADDU.v
// Author        : Cw
// Created On    : 2022-10-17 21:36
// Last Modified : 2022-10-18 19:43
// ---------------------------------------------------------------------------------
// Description   : 
//
//
// -FHDR----------------------------------------------------------------------------
module ysyx_22041752_ADDU (
    input  wire [63: 0] src1,
    input  wire [63: 0] src2,
    output reg  [63: 0] result
);
   
always @(*) begin
    result = src1 + src2;
end

endmodule
