// +FHDR----------------------------------------------------------------------------
//                 Copyright (c) 2022 
//                       ALL RIGHTS RESERVED
// ---------------------------------------------------------------------------------
// Filename      : ysyx_22041752_EXU.v
// Author        : Cw
// Created On    : 2022-11-19 16:16
// Last Modified : 2023-06-02 17:43
// ---------------------------------------------------------------------------------
// Description   : 
//
//
// -FHDR----------------------------------------------------------------------------
`include "ysyx_22041752_mycpu.vh"

module ysyx_22041752_EXU(
    input                                          clk           ,
    input                                          reset         ,

    input                                          ms_allowin    ,
    output                                         es_allowin    ,

    input                                          ds_to_es_valid,
    input  [`ysyx_22041752_DS_TO_ES_BUS_WD -1:0]   ds_to_es_bus  ,

    output                                         es_to_ms_valid,
    output [`ysyx_22041752_ES_TO_MS_BUS_WD -1:0]   es_to_ms_bus  ,

	output [`ysyx_22041752_ES_FORWARD_BUS_WD -1:0] es_forward_bus,

    output                                         data_en       ,
    input                                          data_ready    ,
    output [`ysyx_22041752_SRAM_WEN_WD -1:0]       data_wen      ,
    output [`ysyx_22041752_SRAM_ADDR_WD-1:0]       data_addr     ,
    output [`ysyx_22041752_SRAM_DATA_WD-1:0]       data_wdata    ,

    output                                         flush         ,
    output [`ysyx_22041752_PC_WD-1:0]              flush_pc      ,
    input                                          int_t_i        
);

reg         es_valid      ;
wire        es_ready_go   ;

reg  [`ysyx_22041752_DS_TO_ES_BUS_WD -1:0] ds_to_es_bus_r;  

wire ecall  ;
wire mret   ;
wire mul_u  ;
wire mul_su ;
wire mul_h  ;
wire div_u  ;
wire op_mul ;
wire op_div ;
wire op_rem ;
wire op_add ;
wire op_sub ;
wire op_slt ;
wire op_sltu;
wire op_and ;
wire op_or  ;
wire op_xor ;
wire op_sll ;
wire op_srl ;
wire op_sra ;

wire        res_sext    ;
wire        res_zext    ;
wire        src_shamt   ;
wire        src_pc      ;
wire        src_imm_u   ;
wire        src_4       ;
wire        src_0       ;
wire        src_imm_i   ;
wire        src_imm_s   ;
wire        csrrs       ;
wire        csrrc       ;
wire        src_csr     ;
wire        es_rf_we    ;
wire        es_csr_we   ;
wire        es_mem_we   ;
wire        es_mem_re   ;
wire [ 1:0] es_mem_bytes;
wire [ 5:0] shamt;
wire [19:0] imm_u;
wire [11:0] imm_i;
wire [11:0] imm_s;
wire [11:0] rscsr;
wire [ 4:0] rd;
wire [`ysyx_22041752_RF_DATA_WD-1:0] rs1_value;
wire [`ysyx_22041752_RF_DATA_WD-1:0] rs2_value;
wire [`ysyx_22041752_PC_WD     -1:0] es_pc  ;

assign {ecall         ,
        mret          ,
        div_u         ,
        mul_u         ,
        mul_su        ,
        mul_h         ,
        op_mul        ,
        op_div        ,
        op_rem        ,
        op_add        ,   
        op_sub        ,  
        op_slt        ,  
        op_sltu       ,  
        op_and        ,  
        op_or         ,  
        op_xor        ,  
        op_sll        ,  
        op_srl        ,  
        op_sra        ,  
        res_sext      , 
        res_zext      , 
        shamt         ,  
        src_shamt     ,  
		src_pc        ,	
		src_imm_u     ,  
        src_4         ,  
        src_0         ,  
        src_imm_i     ,  
        src_imm_s     ,  
        src_csr       ,
        rscsr         ,
        es_csr_we     ,
        csrrc         ,
        csrrs         ,
        es_rf_we      ,  
        es_mem_we     ,
        es_mem_re     ,
        es_mem_bytes  ,
        rd            ,  
        imm_s         ,  
        imm_i         ,  
        imm_u         ,  
        rs1_value     ,  
        rs2_value     ,  
        es_pc            
       } = ds_to_es_bus_r;

wire [63:0] alu_src1   ;
wire [63:0] alu_src2   ;
wire [63:0] alu_result ;

assign es_to_ms_bus = {res_sext         ,  
                       res_zext         ,
					   es_mem_bytes     ,  
					   es_mem_re        ,  
					   es_rf_we         ,  
                       rd               ,  
                       alu_result       ,  
                       es_pc               
                      };

reg  [1:0] expfsm_pre;
wire [1:0] expfsm_nxt;
parameter IDLE = 0;
parameter W_MEPC  = 1;
parameter W_MCAUSE= 2;
always @(posedge clk) begin
    if (reset) begin
        expfsm_pre <= IDLE;
    end
    else begin
        expfsm_pre <= expfsm_nxt;
    end
end
assign expfsm_nxt = expfsm_pre == IDLE && (ecall || int_t_o) ? W_MEPC   :
                    expfsm_pre == W_MEPC                     ? W_MCAUSE :
                    expfsm_pre == W_MCAUSE                   ? IDLE     :
                                                               expfsm_pre;

wire mul_out_valid;
wire mul_stall = op_mul && !mul_out_valid && es_valid && !flush;
wire div_out_valid;                                              
wire div_stall = op_rem|op_div && !div_out_valid && es_valid && !flush;
wire mem_stall = data_en && !data_ready;
assign es_ready_go    = expfsm_pre != W_MEPC && !div_stall && !mul_stall && !mem_stall;
assign es_allowin     = !es_valid || es_ready_go && ms_allowin;
assign es_to_ms_valid =  es_valid && es_ready_go &&!flush;
always @(posedge clk) begin
    if (reset) begin
        es_valid <= 1'b0;
    end
    else if (es_allowin) begin
        es_valid <= ds_to_es_valid;
    end
end
always @(posedge clk) begin
    if (reset) begin
        ds_to_es_bus_r <= 0;
    end
    else if(ds_to_es_valid && es_allowin) begin
        ds_to_es_bus_r <= ds_to_es_bus;
    end
end

wire        csr_we   ;
wire [11:0] csr_addr ;
wire [63:0] csr_wdata;
wire [63:0] csr_rdata;
wire        int_t_o  ;

ysyx_22041752_csr U_YSYX_22041752_CSR_0(
    .clk                            ( clk                           ),
    .reset                          ( reset                         ),
    .wen                            ( csr_we                        ),
    .addr                           ( csr_addr                      ),
    .wdata                          ( csr_wdata                     ),
    .rdata                          ( csr_rdata                     ),
    .int_t_i                        ( int_t_i                       ),
    .int_t_o                        ( int_t_o                       )
);
assign csr_we    = es_csr_we || expfsm_pre==W_MEPC || expfsm_pre==W_MCAUSE;
assign csr_addr  = (ecall || int_t_o) && (expfsm_pre==IDLE)    ? `ysyx_22041752_CSR_ADDR_MTVEC  :
                   expfsm_pre==W_MEPC    || mret               ? `ysyx_22041752_CSR_ADDR_MEPC   :
                   expfsm_pre==W_MCAUSE                        ? `ysyx_22041752_CSR_ADDR_MCAUSE :
                                                                 rscsr            ;
assign csr_wdata = expfsm_pre == W_MEPC   ? {32'b0, es_pc} :
                   expfsm_pre == W_MCAUSE ? int_t_o ? 64'h8000_0000_0000_0007: 64'hb :
                   {64{csrrs}} & (rs1_value | csr_rdata) |
                   {64{csrrc}} & (rs1_value &~csr_rdata) |
                   {64{!csrrs && !csrrc}} & rs1_value;

assign flush    = (ecall||mret||int_t_o) && es_valid;
assign flush_pc = csr_rdata[31:0];

assign alu_src1 = src_pc   ? {32'b0, es_pc} : 
                  src_0    ? 64'd0          :
                  res_sext && (op_sll || op_srl || op_sra) ? {32'b0,rs1_value[31:0]} :
                  rs1_value;
  
assign alu_src2 = src_csr   ? csr_rdata :
                  src_4     ? 64'd4 : 
                  src_imm_u ? {{32{imm_u[19]}},imm_u,12'b0} :
                  src_imm_i ? {{52{imm_i[11]}},imm_i} :
                  src_imm_s ? {{52{imm_s[11]}},imm_s} :
                  src_shamt ? {58'b0,shamt} :
                  res_sext && (op_sll || op_srl || op_sra) ? {59'b0,rs2_value[4:0]} :
                  (op_sll || op_srl || op_sra) ? {58'b0,rs2_value[5:0]} :
                  rs2_value;

/* verilator lint_off UNUSEDSIGNAL */
wire [63:0] mem_addr;
/* verilator lint_on UNUSEDSIGNAL */
ysyx_22041752_alu U_ALU_0(
    .clk             ( clk            ),
    .reset           ( reset          ),
    .flush           ( flush          ),
    .mul_u           ( mul_u          ),
    .mul_su          ( mul_su         ),
    .div_u           ( div_u          ),
    .mul_h           ( mul_h          ),
    .op_mul          ( op_mul         ),
    .op_div          ( op_div         ),
    .op_rem          ( op_rem         ),
    .op_add          ( op_add         ),
    .op_sub          ( op_sub         ),
    .op_slt          ( op_slt         ),
    .op_sltu         ( op_sltu        ),
    .op_and          ( op_and         ),
    .op_or           ( op_or          ),
    .op_xor          ( op_xor         ),
    .op_sll          ( op_sll         ),
    .op_srl          ( op_srl         ),
    .op_sra          ( op_sra         ),
    .res_sext        ( res_sext       ),
    .alu_src1        ( alu_src1       ),
    .alu_src2        ( alu_src2       ),
    .alu_result      ( alu_result     ),
    .mem_result      ( mem_addr       ),
    .div_out_valid   ( div_out_valid  ),
    .mul_out_valid   ( mul_out_valid  )
);

assign data_addr= mem_addr[31:0];
assign data_en  = (es_mem_re | es_mem_we) & es_valid;
assign data_wen = es_mem_we && es_valid && es_mem_bytes == 2'b11 ? 8'hff : 
                  es_mem_we && es_valid && es_mem_bytes == 2'b10 ? 8'h0f :
                  es_mem_we && es_valid && es_mem_bytes == 2'b01 ? 8'h03 :
                  es_mem_we && es_valid && es_mem_bytes == 2'b00 ? 8'h01 :
                                                                   8'h00 ;

assign data_wdata = rs2_value;
//forward_bus
wire mem_read_after_write;
wire es_forward_valid;
assign mem_read_after_write = (es_mem_re) && es_valid;
assign es_forward_valid = es_rf_we && es_valid;
assign es_forward_bus = {mem_read_after_write,es_forward_valid,alu_result,rd};

endmodule

